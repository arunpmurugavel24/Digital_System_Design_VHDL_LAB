----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Hian Zing Voon
-- 
-- Create Date: 24.05.2024 11:00:29
-- Design Name: 
-- Module Name: memory_content - Behavioral
-- Project Name: Risc V functional CPU 
-- Description: the functions for Loading the assembler txt file, transforming it into a 
--              32Bit bit_vector and then saving it to the Memory.
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use STD.TEXTIO.ALL;
use WORK.cpu_defs_pack.ALL;
use WORK.mnemonics_pack.ALL;

package mem_defs_pack is  -- Declaration of procedure
procedure filetomemory (
    variable f : in text;
    mem : inout Mem_Type);
end mem_defs_pack;
 
package body mem_defs_pack is -- Content of procedure
procedure filetomemory (
    variable f : in text;
    mem : inout Mem_Type) is 
    variable l : line;
    variable s : string(5 downto 1);  -- The line in the text file MUST be longer than this defined string
    variable int1 : integer; -- bei Read integer, it only takes 1 number, automatically separated by space
    variable int2 : integer; 
    variable int3 : integer;
    variable success : boolean;
          
    begin
        
        -- Read is a 2-step-process; first extract the entire line via "readline", then read part by part via "read"
        while not endfile(f) loop
            readline (f, l);
            success := TRUE;
            
            -- read opcodes
            read(l, s, success);
            
            --read integers after opcodes if they exist
            if success then
                read(l, int1, success);
                if success then
                    read(l, int2, success);
                    if success then
                        read(l, int3, success);
--                        mnemonics_opcode(s);
                        report ("Read line: " & s & "|" & integer'image(int1) & "|" & integer'image(int2) & "|" & integer'image(int3));
                    else 
                        report("Line does not fit the format!");
                    end if;
                end if;
            end if;
---------------------            
--MADE BY Yu-Hung TSAI 
---------------------
        variable Instr_str : string(1 to 32);
        variable opcode_str : string(1 to 7);
        variable rd_str : string(1 to 5);
        variable imm_str : string(1 to 20);        
                                
        if opcode_str = "0110111" then  -- U-type
            imm_str := Instr_str(8 to 32);

            opcode <= bit_vector(opcode_str);
            imm_u <= bit_vector(imm_str);

            binary_instr <= imm_u & rd & opcode;

        elsif opcode_str = "1101111" then  -- J-type
            imm_str := Instr_str(1 to 1) & Instr_str(2 to 10) & Instr_str(11 to 11) & Instr_str(12 to 19) & Instr_str(20 to 31);

            opcode <= bit_vector(opcode_str);
            imm_j <= bit_vector(imm_str);

            binary_instr <= imm_j(20) & imm_j(10 downto 1) & imm_j(11) & imm_j(19 downto 12) & rd & opcode;
        else
            binary_instr <= (others => '0');
        end if;

         
         --------------TEMP-------------------   
--          while not endfile(f) loop
--          readline (f, l);
--          read(l, int1, success);
--          read(l, int2, success);
--          read(l, int3, success);                
--        if success then
--            report ("Read line: " & s & "|" & integer'image(int1) & "|" & integer'image(int2) & "|" & integer'image(int3));
--        else
--            report ("error");
--        end if;

        --------------------------------------
        end loop;
    
--        readline (f, l); 
--        read(l, s, success);
        
--        if success then 
--            report ("---------------!!!!!!!!!-------------" & s);
--        --report("Test");
--        else
--            report ("error");
--        end if; 
        
--        readline (f,l);
--        read(l,s,success);
        
--        if success then
--            report ("scheissssssssssssse" & integer'image(i));
--            report ("---------------!!!----------" & s);
--        else
--            report ("error");
--        end if;
        
--        read(l,i,success);
        
--        if success then
--            report ("kackkkkkkkke" & integer'image(i));
--        else
--            report ("error");
--        end if;
             
end filetomemory;
end mem_defs_pack;

                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        
